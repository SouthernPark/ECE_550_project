module and_32(data_operandA, data_operandB);
	//this module will return the and result of A and B
	input [31:0] data_operandA, data_operandB;


endmodule